* NGSPICE file created from hello_world_hand.ext - technology: sky130A

.subckt hello_world_hand
X0 Y A VGND VSUBS sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=2.4e+06u as=3.25e+11p ps=2.3e+06u w=650000u l=150000u
X1 Y A VPWR NWELL sky130_fd_pr__pfet_01v8 ad=5.5e+11p pd=3.1e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u


