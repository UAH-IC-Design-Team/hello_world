Inverter Simulation
* Include the Sky130 libraries
.lib "/foss/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.include "/foss/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice"


* The following subckt was created by Magic
.subckt hello_world_hand Y A NWELL VSUBS VGND VPWR
X0 Y A VGND VSUBS sky130_fd_pr__nfet_01v8 ad=3.575e+11p pd=2.4e+06u as=3.25e+11p ps=2.3e+06u w=650000u l=150000u
X1 Y A VPWR NWELL sky130_fd_pr__pfet_01v8 ad=5.5e+11p pd=3.1e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
.ends

* instantiate the inverter
Xinv Y A VPWR VGND VGND VPWR hello_world_hand

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
Vin A VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10e-12 2e-09 0e-00

.control
run
set color0 = white
set color1 = black
plot A Y
plot i(Vdd)
.endc

.end
