** sch_path: /foss/designs/hello_world/xschem/hello_world_test.sch
**.subckt hello_world_test
x1 Q VDD VSS Q_n hello_world
V3 VDD GND 1.8V
V4 VSS GND 0
V2 Q GND PULSE 0 1.8V 0 1ns 1ns 10us 20us
**** begin user architecture code
 .lib /foss/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice


.options acct list
.temp 25
*vvcc VDD 0 dc 1.8
*vvss VSS 0 0
.control
*tran 0.1u 60u
dc V2 0 1.8 1m
*plot RST_PLS clk+2 Pulse+4
plot Q Q_n
write hello_world_test.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  hello_world.sym # of pins=4
** sym_path: /foss/designs/hello_world/xschem/hello_world.sym
** sch_path: /foss/designs/hello_world/xschem/hello_world.sch
.subckt hello_world  Q VDD VSS Q_n
*.ipin Q
*.opin Q_n
*.iopin VDD
*.iopin VSS
XM1 Q_n Q VDD VSS sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM2 Q_n Q VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
.ends

.GLOBAL GND
.end
